// transcript from my solution

# NS = red,    EW = red,    time = 0
# NS = red,    EW = green,  time = 75000
# NS = red,    EW = yellow, time = 125000
# NS = red,    EW = red,    time = 145000
# NS = green,  EW = red,    time = 155000
# NS = yellow, EW = red,    time = 205000
# NS = red,    EW = red,    time = 225000
# NS = green,  EW = red,    time = 425000
# NS = yellow, EW = red,    time = 475000
# NS = red,    EW = red,    time = 495000
# NS = red,    EW = green,  time = 505000
# NS = red,    EW = yellow, time = 555000
# NS = red,    EW = red,    time = 575000